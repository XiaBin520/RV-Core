module decoder(
  input         clock,
  input         reset,
  input  [31:0] io_instr,
  output [2:0]  io_immCtrl,
  output [3:0]  io_ctrlModel,
  output [3:0]  io_aluOP,
  output [2:0]  io_aluSrc1Ctrl,
  output [2:0]  io_aluSrc2Ctrl,
  output        io_aluWEn,
  output [2:0]  io_aluWOP,
  output        io_memREn,
  output [2:0]  io_memRCtrl,
  output        io_memWEn,
  output [2:0]  io_memWCtrl,
  output        io_regWEn,
  output [1:0]  io_regWSrc,
  output [4:0]  io_rd,
  output        io_rs1REn,
  output        io_rs2REn,
  output [4:0]  io_rs1,
  output [4:0]  io_rs2
);
  wire [6:0] opcode = io_instr[6:0]; // @[decoder.scala 52:24]
  wire [2:0] funct3 = io_instr[14:12]; // @[decoder.scala 54:24]
  wire [6:0] funct7 = io_instr[31:25]; // @[decoder.scala 57:24]
  wire  _T_3 = 3'h0 == funct3; // @[decoder.scala 125:21]
  wire  _T_4 = 3'h1 == funct3; // @[decoder.scala 125:21]
  wire  _T_5 = 3'h4 == funct3; // @[decoder.scala 125:21]
  wire  _T_6 = 3'h5 == funct3; // @[decoder.scala 125:21]
  wire  _T_7 = 3'h6 == funct3; // @[decoder.scala 125:21]
  wire  _T_8 = 3'h7 == funct3; // @[decoder.scala 125:21]
  wire [3:0] _GEN_0 = 3'h7 == funct3 ? 4'h6 : 4'h0; // @[decoder.scala 125:21 131:33]
  wire [3:0] _GEN_1 = 3'h6 == funct3 ? 4'h5 : _GEN_0; // @[decoder.scala 125:21 130:33]
  wire [3:0] _GEN_2 = 3'h5 == funct3 ? 4'h4 : _GEN_1; // @[decoder.scala 125:21 129:33]
  wire [3:0] _GEN_3 = 3'h4 == funct3 ? 4'h3 : _GEN_2; // @[decoder.scala 125:21 128:33]
  wire [3:0] _GEN_4 = 3'h1 == funct3 ? 4'h2 : _GEN_3; // @[decoder.scala 125:21 127:33]
  wire [3:0] _GEN_5 = 3'h0 == funct3 ? 4'h1 : _GEN_4; // @[decoder.scala 125:21 126:33]
  wire  _T_12 = 3'h2 == funct3; // @[decoder.scala 151:21]
  wire  _T_13 = 3'h3 == funct3; // @[decoder.scala 151:21]
  wire [2:0] _GEN_6 = _T_7 ? 3'h6 : 3'h0; // @[decoder.scala 151:21 158:32]
  wire [2:0] _GEN_7 = _T_6 ? 3'h5 : _GEN_6; // @[decoder.scala 151:21 157:32]
  wire [2:0] _GEN_8 = _T_5 ? 3'h4 : _GEN_7; // @[decoder.scala 151:21 156:32]
  wire [2:0] _GEN_9 = 3'h3 == funct3 ? 3'h7 : _GEN_8; // @[decoder.scala 151:21 155:32]
  wire [2:0] _GEN_10 = 3'h2 == funct3 ? 3'h3 : _GEN_9; // @[decoder.scala 151:21 154:32]
  wire [2:0] _GEN_11 = _T_4 ? 3'h2 : _GEN_10; // @[decoder.scala 151:21 153:32]
  wire [2:0] _GEN_12 = _T_3 ? 3'h1 : _GEN_11; // @[decoder.scala 151:21 152:32]
  wire [2:0] _GEN_13 = _T_13 ? 3'h4 : 3'h0; // @[decoder.scala 173:21 177:32]
  wire [2:0] _GEN_14 = _T_12 ? 3'h3 : _GEN_13; // @[decoder.scala 173:21 176:32]
  wire [2:0] _GEN_15 = _T_4 ? 3'h2 : _GEN_14; // @[decoder.scala 173:21 175:32]
  wire [2:0] _GEN_16 = _T_3 ? 3'h1 : _GEN_15; // @[decoder.scala 173:21 174:32]
  wire [6:0] _T_30 = funct7 & 7'h7e; // @[decoder.scala 206:23]
  wire  _T_31 = 7'h0 == _T_30; // @[decoder.scala 206:23]
  wire [3:0] _GEN_17 = 7'h0 == _T_30 ? 4'h7 : 4'h0; // @[decoder.scala 206:47 207:29]
  wire [3:0] _GEN_18 = 7'h20 == _T_30 ? 4'h9 : 4'h0; // @[decoder.scala 214:52 215:29]
  wire [3:0] _GEN_19 = _T_31 ? 4'h8 : _GEN_18; // @[decoder.scala 211:47 212:29]
  wire [3:0] _GEN_20 = _T_6 ? _GEN_19 : 4'h0; // @[decoder.scala 198:21]
  wire [3:0] _GEN_21 = _T_4 ? _GEN_17 : _GEN_20; // @[decoder.scala 198:21]
  wire [3:0] _GEN_22 = _T_8 ? 4'h6 : _GEN_21; // @[decoder.scala 198:21 204:29]
  wire [3:0] _GEN_23 = _T_7 ? 4'h5 : _GEN_22; // @[decoder.scala 198:21 203:29]
  wire [3:0] _GEN_24 = _T_5 ? 4'h4 : _GEN_23; // @[decoder.scala 198:21 202:29]
  wire [3:0] _GEN_25 = _T_13 ? 4'h3 : _GEN_24; // @[decoder.scala 198:21 201:29]
  wire [3:0] _GEN_26 = _T_12 ? 4'h2 : _GEN_25; // @[decoder.scala 198:21 200:29]
  wire [3:0] _GEN_27 = _T_3 ? 4'h0 : _GEN_26; // @[decoder.scala 198:21 199:29]
  wire [2:0] _GEN_28 = funct7 == 7'h20 ? 3'h5 : 3'h0; // @[decoder.scala 242:46 243:30]
  wire [2:0] _GEN_29 = funct7 == 7'h0 ? 3'h4 : _GEN_28; // @[decoder.scala 239:41 240:30]
  wire [2:0] _GEN_30 = _T_6 ? _GEN_29 : 3'h0; // @[decoder.scala 235:21]
  wire [2:0] _GEN_31 = _T_4 ? 3'h3 : _GEN_30; // @[decoder.scala 235:21 237:30]
  wire [2:0] _GEN_32 = _T_3 ? 3'h1 : _GEN_31; // @[decoder.scala 235:21 236:30]
  wire  _T_44 = 7'h0 == funct7; // @[decoder.scala 268:21]
  wire [3:0] _GEN_35 = _T_6 ? 4'h8 : _GEN_1; // @[decoder.scala 270:25 276:33]
  wire [3:0] _GEN_36 = _T_5 ? 4'h4 : _GEN_35; // @[decoder.scala 270:25 275:33]
  wire [3:0] _GEN_37 = _T_13 ? 4'h3 : _GEN_36; // @[decoder.scala 270:25 274:33]
  wire [3:0] _GEN_38 = _T_12 ? 4'h2 : _GEN_37; // @[decoder.scala 270:25 273:33]
  wire [3:0] _GEN_39 = _T_4 ? 4'h7 : _GEN_38; // @[decoder.scala 270:25 272:33]
  wire [3:0] _GEN_40 = _T_3 ? 4'h0 : _GEN_39; // @[decoder.scala 270:25 271:33]
  wire  _T_53 = 7'h20 == funct7; // @[decoder.scala 268:21]
  wire [3:0] _GEN_41 = _T_6 ? 4'h9 : 4'h0; // @[decoder.scala 282:25 284:33]
  wire [3:0] _GEN_42 = _T_3 ? 4'h1 : _GEN_41; // @[decoder.scala 282:25 283:33]
  wire [3:0] _GEN_43 = 7'h20 == funct7 ? _GEN_42 : 4'h0; // @[decoder.scala 268:21]
  wire [3:0] _GEN_44 = 7'h0 == funct7 ? _GEN_40 : _GEN_43; // @[decoder.scala 268:21]
  wire [2:0] _GEN_45 = _T_53 ? 3'h2 : 3'h0; // @[decoder.scala 305:25 307:38]
  wire [2:0] _GEN_46 = _T_44 ? 3'h1 : _GEN_45; // @[decoder.scala 305:25 306:38]
  wire [2:0] _GEN_47 = _T_44 ? 3'h3 : 3'h0; // @[decoder.scala 311:25 312:38]
  wire [2:0] _GEN_48 = _T_53 ? 3'h5 : 3'h0; // @[decoder.scala 316:25 318:38]
  wire [2:0] _GEN_49 = _T_44 ? 3'h4 : _GEN_48; // @[decoder.scala 316:25 317:38]
  wire [2:0] _GEN_50 = _T_6 ? _GEN_49 : 3'h0; // @[decoder.scala 303:21]
  wire [2:0] _GEN_51 = _T_4 ? _GEN_47 : _GEN_50; // @[decoder.scala 303:21]
  wire [2:0] _GEN_52 = _T_3 ? _GEN_46 : _GEN_51; // @[decoder.scala 303:21]
  wire [2:0] _GEN_53 = 7'h67 == opcode ? 3'h1 : 3'h0; // @[decoder.scala 95:17 339:19]
  wire [3:0] _GEN_54 = 7'h67 == opcode ? 4'h8 : 4'h0; // @[decoder.scala 95:17 340:19]
  wire [1:0] _GEN_56 = 7'h67 == opcode ? 2'h2 : 2'h0; // @[decoder.scala 95:17 342:19]
  wire [2:0] _GEN_57 = 7'h67 == opcode ? 3'h3 : 3'h0; // @[decoder.scala 95:17 343:19]
  wire [1:0] _GEN_59 = 7'h67 == opcode ? 2'h1 : 2'h0; // @[decoder.scala 95:17 345:19]
  wire [2:0] _GEN_60 = 7'h6f == opcode ? 3'h5 : _GEN_53; // @[decoder.scala 95:17 330:19]
  wire [3:0] _GEN_61 = 7'h6f == opcode ? 4'h7 : _GEN_54; // @[decoder.scala 95:17 331:19]
  wire [1:0] _GEN_63 = 7'h6f == opcode ? 2'h2 : _GEN_56; // @[decoder.scala 95:17 333:19]
  wire [2:0] _GEN_64 = 7'h6f == opcode ? 3'h3 : _GEN_57; // @[decoder.scala 95:17 334:19]
  wire  _GEN_65 = 7'h6f == opcode | 7'h67 == opcode; // @[decoder.scala 95:17 335:19]
  wire [1:0] _GEN_66 = 7'h6f == opcode ? 2'h1 : _GEN_59; // @[decoder.scala 95:17 336:19]
  wire [1:0] _GEN_68 = 7'h3b == opcode ? 2'h3 : _GEN_63; // @[decoder.scala 95:17 296:19]
  wire [2:0] _GEN_69 = 7'h3b == opcode ? 3'h2 : _GEN_64; // @[decoder.scala 95:17 297:19]
  wire  _GEN_70 = 7'h3b == opcode | _GEN_65; // @[decoder.scala 298:14 95:17]
  wire [1:0] _GEN_71 = 7'h3b == opcode ? 2'h1 : _GEN_66; // @[decoder.scala 299:15 95:17]
  wire [2:0] _GEN_74 = 7'h3b == opcode ? _GEN_52 : 3'h0; // @[decoder.scala 95:17]
  wire [2:0] _GEN_75 = 7'h3b == opcode ? 3'h0 : _GEN_60; // @[decoder.scala 95:17]
  wire [3:0] _GEN_76 = 7'h3b == opcode ? 4'h0 : _GEN_61; // @[decoder.scala 95:17]
  wire [1:0] _GEN_78 = 7'h33 == opcode ? 2'h3 : _GEN_68; // @[decoder.scala 95:17 262:19]
  wire [2:0] _GEN_79 = 7'h33 == opcode ? 3'h2 : _GEN_69; // @[decoder.scala 95:17 263:19]
  wire  _GEN_80 = 7'h33 == opcode | _GEN_70; // @[decoder.scala 264:14 95:17]
  wire [1:0] _GEN_81 = 7'h33 == opcode ? 2'h1 : _GEN_71; // @[decoder.scala 265:15 95:17]
  wire  _GEN_83 = 7'h33 == opcode | 7'h3b == opcode; // @[decoder.scala 267:14 95:17]
  wire [3:0] _GEN_84 = 7'h33 == opcode ? _GEN_44 : 4'h0; // @[decoder.scala 95:17]
  wire  _GEN_85 = 7'h33 == opcode ? 1'h0 : 7'h3b == opcode; // @[decoder.scala 95:17]
  wire [2:0] _GEN_86 = 7'h33 == opcode ? 3'h0 : _GEN_74; // @[decoder.scala 95:17]
  wire [2:0] _GEN_87 = 7'h33 == opcode ? 3'h0 : _GEN_75; // @[decoder.scala 95:17]
  wire [3:0] _GEN_88 = 7'h33 == opcode ? 4'h0 : _GEN_76; // @[decoder.scala 95:17]
  wire [2:0] _GEN_89 = 7'h1b == opcode ? 3'h1 : _GEN_87; // @[decoder.scala 229:15 95:17]
  wire [1:0] _GEN_90 = 7'h1b == opcode ? 2'h3 : _GEN_78; // @[decoder.scala 95:17 230:19]
  wire [2:0] _GEN_91 = 7'h1b == opcode ? 3'h1 : _GEN_79; // @[decoder.scala 95:17 231:19]
  wire  _GEN_92 = 7'h1b == opcode | _GEN_80; // @[decoder.scala 232:14 95:17]
  wire [1:0] _GEN_93 = 7'h1b == opcode ? 2'h1 : _GEN_81; // @[decoder.scala 233:15 95:17]
  wire [2:0] _GEN_95 = 7'h1b == opcode ? _GEN_32 : _GEN_86; // @[decoder.scala 95:17]
  wire  _GEN_96 = 7'h1b == opcode ? 1'h0 : _GEN_83; // @[decoder.scala 95:17]
  wire [3:0] _GEN_97 = 7'h1b == opcode ? 4'h0 : _GEN_84; // @[decoder.scala 95:17]
  wire  _GEN_98 = 7'h1b == opcode ? 1'h0 : _GEN_85; // @[decoder.scala 95:17]
  wire [3:0] _GEN_99 = 7'h1b == opcode ? 4'h0 : _GEN_88; // @[decoder.scala 95:17]
  wire [2:0] _GEN_100 = 7'h13 == opcode ? 3'h1 : _GEN_89; // @[decoder.scala 95:17 192:19]
  wire [1:0] _GEN_101 = 7'h13 == opcode ? 2'h3 : _GEN_90; // @[decoder.scala 95:17 193:19]
  wire [2:0] _GEN_102 = 7'h13 == opcode ? 3'h1 : _GEN_91; // @[decoder.scala 95:17 194:19]
  wire  _GEN_103 = 7'h13 == opcode | _GEN_92; // @[decoder.scala 95:17 195:19]
  wire [1:0] _GEN_104 = 7'h13 == opcode ? 2'h1 : _GEN_93; // @[decoder.scala 95:17 196:19]
  wire [3:0] _GEN_106 = 7'h13 == opcode ? _GEN_27 : _GEN_97; // @[decoder.scala 95:17]
  wire [2:0] _GEN_107 = 7'h13 == opcode ? 3'h0 : _GEN_95; // @[decoder.scala 95:17]
  wire  _GEN_108 = 7'h13 == opcode ? 1'h0 : _GEN_96; // @[decoder.scala 95:17]
  wire  _GEN_109 = 7'h13 == opcode ? 1'h0 : _GEN_98; // @[decoder.scala 95:17]
  wire [3:0] _GEN_110 = 7'h13 == opcode ? 4'h0 : _GEN_99; // @[decoder.scala 95:17]
  wire [2:0] _GEN_111 = 7'h23 == opcode ? 3'h2 : _GEN_100; // @[decoder.scala 95:17 167:19]
  wire [3:0] _GEN_112 = 7'h23 == opcode ? 4'h0 : _GEN_106; // @[decoder.scala 95:17 168:19]
  wire [1:0] _GEN_113 = 7'h23 == opcode ? 2'h3 : _GEN_101; // @[decoder.scala 95:17 169:19]
  wire [2:0] _GEN_114 = 7'h23 == opcode ? 3'h1 : _GEN_102; // @[decoder.scala 95:17 170:19]
  wire [2:0] _GEN_117 = 7'h23 == opcode ? _GEN_16 : 3'h0; // @[decoder.scala 95:17]
  wire  _GEN_118 = 7'h23 == opcode ? 1'h0 : _GEN_103; // @[decoder.scala 95:17]
  wire [1:0] _GEN_119 = 7'h23 == opcode ? 2'h0 : _GEN_104; // @[decoder.scala 95:17]
  wire [2:0] _GEN_120 = 7'h23 == opcode ? 3'h0 : _GEN_107; // @[decoder.scala 95:17]
  wire  _GEN_121 = 7'h23 == opcode ? 1'h0 : _GEN_108; // @[decoder.scala 95:17]
  wire  _GEN_122 = 7'h23 == opcode ? 1'h0 : _GEN_109; // @[decoder.scala 95:17]
  wire [3:0] _GEN_123 = 7'h23 == opcode ? 4'h0 : _GEN_110; // @[decoder.scala 95:17]
  wire [2:0] _GEN_124 = 7'h3 == opcode ? 3'h1 : _GEN_111; // @[decoder.scala 95:17 143:19]
  wire [3:0] _GEN_125 = 7'h3 == opcode ? 4'h0 : _GEN_112; // @[decoder.scala 95:17 144:19]
  wire [1:0] _GEN_126 = 7'h3 == opcode ? 2'h3 : _GEN_113; // @[decoder.scala 95:17 145:19]
  wire [2:0] _GEN_127 = 7'h3 == opcode ? 3'h1 : _GEN_114; // @[decoder.scala 95:17 146:19]
  wire  _GEN_129 = 7'h3 == opcode | _GEN_118; // @[decoder.scala 95:17 148:19]
  wire [1:0] _GEN_130 = 7'h3 == opcode ? 2'h2 : _GEN_119; // @[decoder.scala 95:17 149:19]
  wire [2:0] _GEN_132 = 7'h3 == opcode ? _GEN_12 : 3'h0; // @[decoder.scala 95:17]
  wire  _GEN_133 = 7'h3 == opcode ? 1'h0 : 7'h23 == opcode; // @[decoder.scala 95:17]
  wire [2:0] _GEN_134 = 7'h3 == opcode ? 3'h0 : _GEN_117; // @[decoder.scala 95:17]
  wire [2:0] _GEN_135 = 7'h3 == opcode ? 3'h0 : _GEN_120; // @[decoder.scala 95:17]
  wire  _GEN_136 = 7'h3 == opcode ? 1'h0 : _GEN_121; // @[decoder.scala 95:17]
  wire  _GEN_137 = 7'h3 == opcode ? 1'h0 : _GEN_122; // @[decoder.scala 95:17]
  wire [3:0] _GEN_138 = 7'h3 == opcode ? 4'h0 : _GEN_123; // @[decoder.scala 95:17]
  wire [2:0] _GEN_139 = 7'h63 == opcode ? 3'h3 : _GEN_124; // @[decoder.scala 122:15 95:17]
  wire  _GEN_141 = 7'h63 == opcode | _GEN_136; // @[decoder.scala 124:15 95:17]
  wire [3:0] _GEN_142 = 7'h63 == opcode ? _GEN_5 : _GEN_138; // @[decoder.scala 95:17]
  wire [3:0] _GEN_143 = 7'h63 == opcode ? 4'h0 : _GEN_125; // @[decoder.scala 95:17]
  wire [1:0] _GEN_144 = 7'h63 == opcode ? 2'h0 : _GEN_126; // @[decoder.scala 95:17]
  wire [2:0] _GEN_145 = 7'h63 == opcode ? 3'h0 : _GEN_127; // @[decoder.scala 95:17]
  wire  _GEN_146 = 7'h63 == opcode ? 1'h0 : 7'h3 == opcode; // @[decoder.scala 95:17]
  wire  _GEN_147 = 7'h63 == opcode ? 1'h0 : _GEN_129; // @[decoder.scala 95:17]
  wire [1:0] _GEN_148 = 7'h63 == opcode ? 2'h0 : _GEN_130; // @[decoder.scala 95:17]
  wire [2:0] _GEN_149 = 7'h63 == opcode ? 3'h0 : _GEN_132; // @[decoder.scala 95:17]
  wire  _GEN_150 = 7'h63 == opcode ? 1'h0 : _GEN_133; // @[decoder.scala 95:17]
  wire [2:0] _GEN_151 = 7'h63 == opcode ? 3'h0 : _GEN_134; // @[decoder.scala 95:17]
  wire [2:0] _GEN_152 = 7'h63 == opcode ? 3'h0 : _GEN_135; // @[decoder.scala 95:17]
  wire  _GEN_153 = 7'h63 == opcode ? 1'h0 : _GEN_137; // @[decoder.scala 95:17]
  wire [2:0] _GEN_154 = 7'h17 == opcode ? 3'h4 : _GEN_139; // @[decoder.scala 95:17 107:19]
  wire [3:0] _GEN_155 = 7'h17 == opcode ? 4'h0 : _GEN_143; // @[decoder.scala 95:17 108:19]
  wire [1:0] _GEN_156 = 7'h17 == opcode ? 2'h2 : _GEN_144; // @[decoder.scala 95:17 109:19]
  wire [2:0] _GEN_157 = 7'h17 == opcode ? 3'h1 : _GEN_145; // @[decoder.scala 95:17 110:19]
  wire  _GEN_158 = 7'h17 == opcode | _GEN_147; // @[decoder.scala 95:17 111:19]
  wire [1:0] _GEN_159 = 7'h17 == opcode ? 2'h1 : _GEN_148; // @[decoder.scala 95:17 112:19]
  wire  _GEN_161 = 7'h17 == opcode ? 1'h0 : _GEN_141; // @[decoder.scala 95:17]
  wire [3:0] _GEN_162 = 7'h17 == opcode ? 4'h0 : _GEN_142; // @[decoder.scala 95:17]
  wire  _GEN_163 = 7'h17 == opcode ? 1'h0 : _GEN_146; // @[decoder.scala 95:17]
  wire [2:0] _GEN_164 = 7'h17 == opcode ? 3'h0 : _GEN_149; // @[decoder.scala 95:17]
  wire  _GEN_165 = 7'h17 == opcode ? 1'h0 : _GEN_150; // @[decoder.scala 95:17]
  wire [2:0] _GEN_166 = 7'h17 == opcode ? 3'h0 : _GEN_151; // @[decoder.scala 95:17]
  wire [2:0] _GEN_167 = 7'h17 == opcode ? 3'h0 : _GEN_152; // @[decoder.scala 95:17]
  wire  _GEN_168 = 7'h17 == opcode ? 1'h0 : _GEN_153; // @[decoder.scala 95:17]
  wire [1:0] aluSrc1Ctrl = 7'h37 == opcode ? 2'h1 : _GEN_156; // @[decoder.scala 95:17 100:19]
  assign io_immCtrl = 7'h37 == opcode ? 3'h4 : _GEN_154; // @[decoder.scala 95:17 98:19]
  assign io_ctrlModel = 7'h37 == opcode ? 4'h0 : _GEN_162; // @[decoder.scala 95:17]
  assign io_aluOP = 7'h37 == opcode ? 4'h0 : _GEN_155; // @[decoder.scala 95:17 99:19]
  assign io_aluSrc1Ctrl = {{1'd0}, aluSrc1Ctrl}; // @[decoder.scala 402:20]
  assign io_aluSrc2Ctrl = 7'h37 == opcode ? 3'h1 : _GEN_157; // @[decoder.scala 95:17 101:19]
  assign io_aluWEn = 7'h37 == opcode ? 1'h0 : _GEN_168; // @[decoder.scala 95:17]
  assign io_aluWOP = 7'h37 == opcode ? 3'h0 : _GEN_167; // @[decoder.scala 95:17]
  assign io_memREn = 7'h37 == opcode ? 1'h0 : _GEN_163; // @[decoder.scala 95:17]
  assign io_memRCtrl = 7'h37 == opcode ? 3'h0 : _GEN_164; // @[decoder.scala 95:17]
  assign io_memWEn = 7'h37 == opcode ? 1'h0 : _GEN_165; // @[decoder.scala 95:17]
  assign io_memWCtrl = 7'h37 == opcode ? 3'h0 : _GEN_166; // @[decoder.scala 95:17]
  assign io_regWEn = 7'h37 == opcode | _GEN_158; // @[decoder.scala 95:17 102:19]
  assign io_regWSrc = 7'h37 == opcode ? 2'h1 : _GEN_159; // @[decoder.scala 95:17 103:19]
  assign io_rd = io_instr[11:7]; // @[decoder.scala 53:24]
  assign io_rs1REn = 7'h37 == opcode ? 1'h0 : _GEN_161; // @[decoder.scala 95:17]
  assign io_rs2REn = 7'h37 == opcode ? 1'h0 : _GEN_161; // @[decoder.scala 95:17]
  assign io_rs1 = io_instr[19:15]; // @[decoder.scala 55:24]
  assign io_rs2 = io_instr[24:20]; // @[decoder.scala 56:24]
endmodule
