module Decoder(
  input  [31:0] io_INSTRIN_Instr,
  output [2:0]  io_IMMCTRL_ImmCtrl,
  output [3:0]  io_JUMPCTRL_JumpCtrl,
  output [3:0]  io_ALUCTRL_ALUOP,
  output [2:0]  io_ALUCTRL_ALUData1Ctrl,
  output [2:0]  io_ALUCTRL_ALUData2Ctrl,
  output        io_ALUCTRL_WordALUEn,
  output [2:0]  io_ALUCTRL_WordALUOP,
  output        io_MEMCTRL_REn,
  output [2:0]  io_MEMCTRL_RCtrl,
  output        io_MEMCTRL_WEn,
  output [2:0]  io_MEMCTRL_WCtrl,
  output        io_REGWRITE_WEn,
  output [4:0]  io_REGWRITE_Rd,
  output [4:0]  io_REGREAD_A_Rs1,
  output [4:0]  io_REGREAD_A_Rs2,
  output        io_REGREAD_B_Rs1En,
  output        io_REGREAD_B_Rs2En
);
  wire [6:0] Opcode = io_INSTRIN_Instr[6:0]; // @[Decoder.scala 93:32]
  wire [2:0] Funct3 = io_INSTRIN_Instr[14:12]; // @[Decoder.scala 95:32]
  wire [6:0] Funct7 = io_INSTRIN_Instr[31:25]; // @[Decoder.scala 98:32]
  wire  _T_3 = 3'h0 == Funct3; // @[Decoder.scala 161:21]
  wire  _T_4 = 3'h1 == Funct3; // @[Decoder.scala 161:21]
  wire  _T_5 = 3'h4 == Funct3; // @[Decoder.scala 161:21]
  wire  _T_6 = 3'h5 == Funct3; // @[Decoder.scala 161:21]
  wire  _T_7 = 3'h6 == Funct3; // @[Decoder.scala 161:21]
  wire  _T_8 = 3'h7 == Funct3; // @[Decoder.scala 161:21]
  wire [3:0] _GEN_0 = 3'h7 == Funct3 ? 4'h6 : 4'h0; // @[Decoder.scala 161:21 167:32]
  wire [3:0] _GEN_1 = 3'h6 == Funct3 ? 4'h5 : _GEN_0; // @[Decoder.scala 161:21 166:32]
  wire [3:0] _GEN_2 = 3'h5 == Funct3 ? 4'h4 : _GEN_1; // @[Decoder.scala 161:21 165:32]
  wire [3:0] _GEN_3 = 3'h4 == Funct3 ? 4'h3 : _GEN_2; // @[Decoder.scala 161:21 164:32]
  wire [3:0] _GEN_4 = 3'h1 == Funct3 ? 4'h2 : _GEN_3; // @[Decoder.scala 161:21 163:32]
  wire [3:0] _GEN_5 = 3'h0 == Funct3 ? 4'h1 : _GEN_4; // @[Decoder.scala 161:21 162:32]
  wire  _T_12 = 3'h2 == Funct3; // @[Decoder.scala 186:21]
  wire  _T_13 = 3'h3 == Funct3; // @[Decoder.scala 186:21]
  wire [2:0] _GEN_6 = _T_7 ? 3'h6 : 3'h0; // @[Decoder.scala 186:21 193:32]
  wire [2:0] _GEN_7 = _T_6 ? 3'h5 : _GEN_6; // @[Decoder.scala 186:21 192:32]
  wire [2:0] _GEN_8 = _T_5 ? 3'h4 : _GEN_7; // @[Decoder.scala 186:21 191:32]
  wire [2:0] _GEN_9 = 3'h3 == Funct3 ? 3'h7 : _GEN_8; // @[Decoder.scala 186:21 190:32]
  wire [2:0] _GEN_10 = 3'h2 == Funct3 ? 3'h3 : _GEN_9; // @[Decoder.scala 186:21 189:32]
  wire [2:0] _GEN_11 = _T_4 ? 3'h2 : _GEN_10; // @[Decoder.scala 186:21 188:32]
  wire [2:0] _GEN_12 = _T_3 ? 3'h1 : _GEN_11; // @[Decoder.scala 186:21 187:32]
  wire [2:0] _GEN_13 = _T_13 ? 3'h4 : 3'h0; // @[Decoder.scala 209:21 213:32]
  wire [2:0] _GEN_14 = _T_12 ? 3'h3 : _GEN_13; // @[Decoder.scala 209:21 212:32]
  wire [2:0] _GEN_15 = _T_4 ? 3'h2 : _GEN_14; // @[Decoder.scala 209:21 211:32]
  wire [2:0] _GEN_16 = _T_3 ? 3'h1 : _GEN_15; // @[Decoder.scala 209:21 210:32]
  wire [6:0] _T_30 = Funct7 & 7'h7e; // @[Decoder.scala 240:36]
  wire  _T_31 = 7'h0 == _T_30; // @[Decoder.scala 240:36]
  wire [3:0] _GEN_17 = 7'h0 == _T_30 ? 4'h7 : 4'h0; // @[Decoder.scala 240:{60,67}]
  wire [3:0] _GEN_18 = 7'h20 == _T_30 ? 4'h9 : 4'h0; // @[Decoder.scala 242:{60,67}]
  wire [3:0] _GEN_19 = _T_31 ? 4'h8 : _GEN_18; // @[Decoder.scala 241:{60,67}]
  wire [3:0] _GEN_20 = _T_6 ? _GEN_19 : 4'h0; // @[Decoder.scala 233:21]
  wire [3:0] _GEN_21 = _T_4 ? _GEN_17 : _GEN_20; // @[Decoder.scala 233:21]
  wire [3:0] _GEN_22 = _T_8 ? 4'h6 : _GEN_21; // @[Decoder.scala 233:21 239:29]
  wire [3:0] _GEN_23 = _T_7 ? 4'h5 : _GEN_22; // @[Decoder.scala 233:21 238:29]
  wire [3:0] _GEN_24 = _T_5 ? 4'h4 : _GEN_23; // @[Decoder.scala 233:21 237:29]
  wire [3:0] _GEN_25 = _T_13 ? 4'h3 : _GEN_24; // @[Decoder.scala 233:21 236:29]
  wire [3:0] _GEN_26 = _T_12 ? 4'h2 : _GEN_25; // @[Decoder.scala 233:21 235:29]
  wire [3:0] _GEN_27 = _T_3 ? 4'h0 : _GEN_26; // @[Decoder.scala 233:21 234:29]
  wire [2:0] _GEN_28 = Funct7 == 7'h20 ? 3'h5 : 3'h0; // @[Decoder.scala 263:{53,64}]
  wire [2:0] _GEN_29 = Funct7 == 7'h0 ? 3'h4 : _GEN_28; // @[Decoder.scala 262:{53,64}]
  wire [2:0] _GEN_30 = _T_6 ? _GEN_29 : 3'h0; // @[Decoder.scala 259:21]
  wire [2:0] _GEN_31 = _T_4 ? 3'h3 : _GEN_30; // @[Decoder.scala 259:21 261:33]
  wire [2:0] _GEN_32 = _T_3 ? 3'h1 : _GEN_31; // @[Decoder.scala 259:21 260:33]
  wire  _T_44 = 7'h0 == Funct7; // @[Decoder.scala 285:21]
  wire [3:0] _GEN_35 = _T_6 ? 4'h8 : _GEN_1; // @[Decoder.scala 287:25 293:33]
  wire [3:0] _GEN_36 = _T_5 ? 4'h4 : _GEN_35; // @[Decoder.scala 287:25 292:33]
  wire [3:0] _GEN_37 = _T_13 ? 4'h3 : _GEN_36; // @[Decoder.scala 287:25 291:33]
  wire [3:0] _GEN_38 = _T_12 ? 4'h2 : _GEN_37; // @[Decoder.scala 287:25 290:33]
  wire [3:0] _GEN_39 = _T_4 ? 4'h7 : _GEN_38; // @[Decoder.scala 287:25 289:33]
  wire [3:0] _GEN_40 = _T_3 ? 4'h0 : _GEN_39; // @[Decoder.scala 287:25 288:33]
  wire  _T_53 = 7'h20 == Funct7; // @[Decoder.scala 285:21]
  wire [3:0] _GEN_41 = _T_6 ? 4'h9 : 4'h0; // @[Decoder.scala 299:25 301:33]
  wire [3:0] _GEN_42 = _T_3 ? 4'h1 : _GEN_41; // @[Decoder.scala 299:25 300:33]
  wire [3:0] _GEN_43 = 7'h20 == Funct7 ? _GEN_42 : 4'h0; // @[Decoder.scala 285:21]
  wire [3:0] _GEN_44 = 7'h0 == Funct7 ? _GEN_40 : _GEN_43; // @[Decoder.scala 285:21]
  wire [2:0] _GEN_45 = _T_53 ? 3'h2 : 3'h0; // @[Decoder.scala 321:25 323:41]
  wire [2:0] _GEN_46 = _T_44 ? 3'h1 : _GEN_45; // @[Decoder.scala 321:25 322:41]
  wire [2:0] _GEN_47 = _T_44 ? 3'h3 : 3'h0; // @[Decoder.scala 327:25 328:41]
  wire [2:0] _GEN_48 = _T_53 ? 3'h5 : 3'h0; // @[Decoder.scala 332:25 334:41]
  wire [2:0] _GEN_49 = _T_44 ? 3'h4 : _GEN_48; // @[Decoder.scala 332:25 333:41]
  wire [2:0] _GEN_50 = _T_6 ? _GEN_49 : 3'h0; // @[Decoder.scala 319:21]
  wire [2:0] _GEN_51 = _T_4 ? _GEN_47 : _GEN_50; // @[Decoder.scala 319:21]
  wire [2:0] _GEN_52 = _T_3 ? _GEN_46 : _GEN_51; // @[Decoder.scala 319:21]
  wire [2:0] _GEN_53 = 7'h67 == Opcode ? 3'h1 : 3'h0; // @[Decoder.scala 133:17 354:19]
  wire [3:0] _GEN_54 = 7'h67 == Opcode ? 4'h8 : 4'h0; // @[Decoder.scala 133:17 355:19]
  wire [1:0] _GEN_56 = 7'h67 == Opcode ? 2'h2 : 2'h0; // @[Decoder.scala 133:17 357:20]
  wire [2:0] _GEN_57 = 7'h67 == Opcode ? 3'h3 : 3'h0; // @[Decoder.scala 133:17 358:20]
  wire [2:0] _GEN_59 = 7'h6f == Opcode ? 3'h5 : _GEN_53; // @[Decoder.scala 133:17 346:19]
  wire [3:0] _GEN_60 = 7'h6f == Opcode ? 4'h7 : _GEN_54; // @[Decoder.scala 133:17 347:19]
  wire [1:0] _GEN_62 = 7'h6f == Opcode ? 2'h2 : _GEN_56; // @[Decoder.scala 133:17 349:20]
  wire [2:0] _GEN_63 = 7'h6f == Opcode ? 3'h3 : _GEN_57; // @[Decoder.scala 133:17 350:20]
  wire  _GEN_64 = 7'h6f == Opcode | 7'h67 == Opcode; // @[Decoder.scala 133:17 351:14]
  wire  _GEN_65 = 7'h6f == Opcode ? 1'h0 : 7'h67 == Opcode; // @[Decoder.scala 133:17]
  wire [1:0] _GEN_66 = 7'h3b == Opcode ? 2'h3 : _GEN_62; // @[Decoder.scala 133:17 313:20]
  wire [2:0] _GEN_67 = 7'h3b == Opcode ? 3'h2 : _GEN_63; // @[Decoder.scala 133:17 314:20]
  wire  _GEN_68 = 7'h3b == Opcode | _GEN_64; // @[Decoder.scala 133:17 315:14]
  wire  _GEN_69 = 7'h3b == Opcode | _GEN_65; // @[Decoder.scala 133:17 316:14]
  wire [2:0] _GEN_71 = 7'h3b == Opcode ? _GEN_52 : 3'h0; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_72 = 7'h3b == Opcode ? 3'h0 : _GEN_59; // @[Decoder.scala 133:17]
  wire [3:0] _GEN_73 = 7'h3b == Opcode ? 4'h0 : _GEN_60; // @[Decoder.scala 133:17]
  wire [1:0] _GEN_75 = 7'h33 == Opcode ? 2'h3 : _GEN_66; // @[Decoder.scala 133:17 280:20]
  wire [2:0] _GEN_76 = 7'h33 == Opcode ? 3'h2 : _GEN_67; // @[Decoder.scala 133:17 281:20]
  wire  _GEN_77 = 7'h33 == Opcode | _GEN_68; // @[Decoder.scala 133:17 282:14]
  wire  _GEN_78 = 7'h33 == Opcode | _GEN_69; // @[Decoder.scala 133:17 283:14]
  wire  _GEN_79 = 7'h33 == Opcode | 7'h3b == Opcode; // @[Decoder.scala 133:17 284:14]
  wire [3:0] _GEN_80 = 7'h33 == Opcode ? _GEN_44 : 4'h0; // @[Decoder.scala 133:17]
  wire  _GEN_81 = 7'h33 == Opcode ? 1'h0 : 7'h3b == Opcode; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_82 = 7'h33 == Opcode ? 3'h0 : _GEN_71; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_83 = 7'h33 == Opcode ? 3'h0 : _GEN_72; // @[Decoder.scala 133:17]
  wire [3:0] _GEN_84 = 7'h33 == Opcode ? 4'h0 : _GEN_73; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_85 = 7'h1b == Opcode ? 3'h1 : _GEN_83; // @[Decoder.scala 133:17 253:19]
  wire [1:0] _GEN_86 = 7'h1b == Opcode ? 2'h3 : _GEN_75; // @[Decoder.scala 133:17 254:20]
  wire [2:0] _GEN_87 = 7'h1b == Opcode ? 3'h1 : _GEN_76; // @[Decoder.scala 133:17 255:20]
  wire  _GEN_88 = 7'h1b == Opcode | _GEN_77; // @[Decoder.scala 133:17 256:17]
  wire  _GEN_89 = 7'h1b == Opcode | _GEN_78; // @[Decoder.scala 133:17 257:17]
  wire  _GEN_90 = 7'h1b == Opcode | _GEN_81; // @[Decoder.scala 133:17 258:17]
  wire [2:0] _GEN_91 = 7'h1b == Opcode ? _GEN_32 : _GEN_82; // @[Decoder.scala 133:17]
  wire  _GEN_92 = 7'h1b == Opcode ? 1'h0 : _GEN_79; // @[Decoder.scala 133:17]
  wire [3:0] _GEN_93 = 7'h1b == Opcode ? 4'h0 : _GEN_80; // @[Decoder.scala 133:17]
  wire [3:0] _GEN_94 = 7'h1b == Opcode ? 4'h0 : _GEN_84; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_95 = 7'h13 == Opcode ? 3'h1 : _GEN_85; // @[Decoder.scala 133:17 228:19]
  wire [1:0] _GEN_96 = 7'h13 == Opcode ? 2'h3 : _GEN_86; // @[Decoder.scala 133:17 229:20]
  wire [2:0] _GEN_97 = 7'h13 == Opcode ? 3'h1 : _GEN_87; // @[Decoder.scala 133:17 230:20]
  wire  _GEN_98 = 7'h13 == Opcode | _GEN_88; // @[Decoder.scala 133:17 231:14]
  wire  _GEN_99 = 7'h13 == Opcode | _GEN_89; // @[Decoder.scala 133:17 232:14]
  wire [3:0] _GEN_100 = 7'h13 == Opcode ? _GEN_27 : _GEN_93; // @[Decoder.scala 133:17]
  wire  _GEN_101 = 7'h13 == Opcode ? 1'h0 : _GEN_90; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_102 = 7'h13 == Opcode ? 3'h0 : _GEN_91; // @[Decoder.scala 133:17]
  wire  _GEN_103 = 7'h13 == Opcode ? 1'h0 : _GEN_92; // @[Decoder.scala 133:17]
  wire [3:0] _GEN_104 = 7'h13 == Opcode ? 4'h0 : _GEN_94; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_105 = 7'h23 == Opcode ? 3'h2 : _GEN_95; // @[Decoder.scala 133:17 202:19]
  wire [3:0] _GEN_106 = 7'h23 == Opcode ? 4'h0 : _GEN_100; // @[Decoder.scala 133:17 203:20]
  wire [1:0] _GEN_107 = 7'h23 == Opcode ? 2'h3 : _GEN_96; // @[Decoder.scala 133:17 204:20]
  wire [2:0] _GEN_108 = 7'h23 == Opcode ? 3'h1 : _GEN_97; // @[Decoder.scala 133:17 205:20]
  wire  _GEN_110 = 7'h23 == Opcode | _GEN_99; // @[Decoder.scala 133:17 207:14]
  wire  _GEN_111 = 7'h23 == Opcode | _GEN_103; // @[Decoder.scala 133:17 208:14]
  wire [2:0] _GEN_112 = 7'h23 == Opcode ? _GEN_16 : 3'h0; // @[Decoder.scala 133:17]
  wire  _GEN_113 = 7'h23 == Opcode ? 1'h0 : _GEN_98; // @[Decoder.scala 133:17]
  wire  _GEN_114 = 7'h23 == Opcode ? 1'h0 : _GEN_101; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_115 = 7'h23 == Opcode ? 3'h0 : _GEN_102; // @[Decoder.scala 133:17]
  wire [3:0] _GEN_116 = 7'h23 == Opcode ? 4'h0 : _GEN_104; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_117 = 7'h3 == Opcode ? 3'h1 : _GEN_105; // @[Decoder.scala 133:17 179:19]
  wire [3:0] _GEN_118 = 7'h3 == Opcode ? 4'h0 : _GEN_106; // @[Decoder.scala 133:17 180:19]
  wire [1:0] _GEN_119 = 7'h3 == Opcode ? 2'h3 : _GEN_107; // @[Decoder.scala 133:17 181:20]
  wire [2:0] _GEN_120 = 7'h3 == Opcode ? 3'h1 : _GEN_108; // @[Decoder.scala 133:17 182:20]
  wire  _GEN_122 = 7'h3 == Opcode | _GEN_113; // @[Decoder.scala 133:17 184:14]
  wire  _GEN_123 = 7'h3 == Opcode | _GEN_110; // @[Decoder.scala 133:17 185:14]
  wire [2:0] _GEN_124 = 7'h3 == Opcode ? _GEN_12 : 3'h0; // @[Decoder.scala 133:17]
  wire  _GEN_125 = 7'h3 == Opcode ? 1'h0 : 7'h23 == Opcode; // @[Decoder.scala 133:17]
  wire  _GEN_126 = 7'h3 == Opcode ? 1'h0 : _GEN_111; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_127 = 7'h3 == Opcode ? 3'h0 : _GEN_112; // @[Decoder.scala 133:17]
  wire  _GEN_128 = 7'h3 == Opcode ? 1'h0 : _GEN_114; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_129 = 7'h3 == Opcode ? 3'h0 : _GEN_115; // @[Decoder.scala 133:17]
  wire [3:0] _GEN_130 = 7'h3 == Opcode ? 4'h0 : _GEN_116; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_131 = 7'h63 == Opcode ? 3'h3 : _GEN_117; // @[Decoder.scala 133:17 158:15]
  wire  _GEN_132 = 7'h63 == Opcode | _GEN_123; // @[Decoder.scala 133:17 159:15]
  wire  _GEN_133 = 7'h63 == Opcode | _GEN_126; // @[Decoder.scala 133:17 160:15]
  wire [3:0] _GEN_134 = 7'h63 == Opcode ? _GEN_5 : _GEN_130; // @[Decoder.scala 133:17]
  wire [3:0] _GEN_135 = 7'h63 == Opcode ? 4'h0 : _GEN_118; // @[Decoder.scala 133:17]
  wire [1:0] _GEN_136 = 7'h63 == Opcode ? 2'h0 : _GEN_119; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_137 = 7'h63 == Opcode ? 3'h0 : _GEN_120; // @[Decoder.scala 133:17]
  wire  _GEN_138 = 7'h63 == Opcode ? 1'h0 : 7'h3 == Opcode; // @[Decoder.scala 133:17]
  wire  _GEN_139 = 7'h63 == Opcode ? 1'h0 : _GEN_122; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_140 = 7'h63 == Opcode ? 3'h0 : _GEN_124; // @[Decoder.scala 133:17]
  wire  _GEN_141 = 7'h63 == Opcode ? 1'h0 : _GEN_125; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_142 = 7'h63 == Opcode ? 3'h0 : _GEN_127; // @[Decoder.scala 133:17]
  wire  _GEN_143 = 7'h63 == Opcode ? 1'h0 : _GEN_128; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_144 = 7'h63 == Opcode ? 3'h0 : _GEN_129; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_145 = 7'h17 == Opcode ? 3'h4 : _GEN_131; // @[Decoder.scala 133:17 144:19]
  wire [3:0] _GEN_146 = 7'h17 == Opcode ? 4'h0 : _GEN_135; // @[Decoder.scala 133:17 145:19]
  wire [1:0] _GEN_147 = 7'h17 == Opcode ? 2'h2 : _GEN_136; // @[Decoder.scala 133:17 146:20]
  wire [2:0] _GEN_148 = 7'h17 == Opcode ? 3'h1 : _GEN_137; // @[Decoder.scala 133:17 147:20]
  wire  _GEN_149 = 7'h17 == Opcode | _GEN_139; // @[Decoder.scala 133:17 148:19]
  wire  _GEN_150 = 7'h17 == Opcode ? 1'h0 : _GEN_132; // @[Decoder.scala 133:17]
  wire  _GEN_151 = 7'h17 == Opcode ? 1'h0 : _GEN_133; // @[Decoder.scala 133:17]
  wire [3:0] _GEN_152 = 7'h17 == Opcode ? 4'h0 : _GEN_134; // @[Decoder.scala 133:17]
  wire  _GEN_153 = 7'h17 == Opcode ? 1'h0 : _GEN_138; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_154 = 7'h17 == Opcode ? 3'h0 : _GEN_140; // @[Decoder.scala 133:17]
  wire  _GEN_155 = 7'h17 == Opcode ? 1'h0 : _GEN_141; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_156 = 7'h17 == Opcode ? 3'h0 : _GEN_142; // @[Decoder.scala 133:17]
  wire  _GEN_157 = 7'h17 == Opcode ? 1'h0 : _GEN_143; // @[Decoder.scala 133:17]
  wire [2:0] _GEN_158 = 7'h17 == Opcode ? 3'h0 : _GEN_144; // @[Decoder.scala 133:17]
  wire [1:0] ALUData1Ctrl = 7'h37 == Opcode ? 2'h1 : _GEN_147; // @[Decoder.scala 133:17 138:20]
  assign io_IMMCTRL_ImmCtrl = 7'h37 == Opcode ? 3'h4 : _GEN_145; // @[Decoder.scala 133:17 136:20]
  assign io_JUMPCTRL_JumpCtrl = 7'h37 == Opcode ? 4'h0 : _GEN_152; // @[Decoder.scala 133:17]
  assign io_ALUCTRL_ALUOP = 7'h37 == Opcode ? 4'h0 : _GEN_146; // @[Decoder.scala 133:17 137:20]
  assign io_ALUCTRL_ALUData1Ctrl = {{1'd0}, ALUData1Ctrl}; // @[Decoder.scala 419:27]
  assign io_ALUCTRL_ALUData2Ctrl = 7'h37 == Opcode ? 3'h1 : _GEN_148; // @[Decoder.scala 133:17 139:20]
  assign io_ALUCTRL_WordALUEn = 7'h37 == Opcode ? 1'h0 : _GEN_157; // @[Decoder.scala 133:17]
  assign io_ALUCTRL_WordALUOP = 7'h37 == Opcode ? 3'h0 : _GEN_158; // @[Decoder.scala 133:17]
  assign io_MEMCTRL_REn = 7'h37 == Opcode ? 1'h0 : _GEN_153; // @[Decoder.scala 133:17]
  assign io_MEMCTRL_RCtrl = 7'h37 == Opcode ? 3'h0 : _GEN_154; // @[Decoder.scala 133:17]
  assign io_MEMCTRL_WEn = 7'h37 == Opcode ? 1'h0 : _GEN_155; // @[Decoder.scala 133:17]
  assign io_MEMCTRL_WCtrl = 7'h37 == Opcode ? 3'h0 : _GEN_156; // @[Decoder.scala 133:17]
  assign io_REGWRITE_WEn = 7'h37 == Opcode | _GEN_149; // @[Decoder.scala 133:17 140:20]
  assign io_REGWRITE_Rd = io_INSTRIN_Instr[11:7]; // @[Decoder.scala 94:32]
  assign io_REGREAD_A_Rs1 = io_INSTRIN_Instr[19:15]; // @[Decoder.scala 96:32]
  assign io_REGREAD_A_Rs2 = io_INSTRIN_Instr[24:20]; // @[Decoder.scala 97:32]
  assign io_REGREAD_B_Rs1En = 7'h37 == Opcode ? 1'h0 : _GEN_150; // @[Decoder.scala 133:17]
  assign io_REGREAD_B_Rs2En = 7'h37 == Opcode ? 1'h0 : _GEN_151; // @[Decoder.scala 133:17]
endmodule
